library ieee;
use ieee.std_logic_1164.all;

entity div6_e is
port(
		en_i: in std_logic;
		clk_i: in std_logic;
		rb_i: in std_logic;
		c_o: out std_logic
	);
end div6_e;
