library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity div25meg_e is
  port (
    clk_i : in     std_logic;
    div_o : out    std_logic;
    rb_i  : in     std_logic);
end entity div25meg_e;



