library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity div4_e is
port(
		en_i: IN std_logic;
		clk_i: IN std_logic;
		rb_i: IN std_logic;
		c_o: OUT std_logic
	);
end div4_e;
