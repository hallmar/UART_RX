library IEEE;
    use IEEE.STD_LOGIC_1164.all;
use ieee.numeric_std.all;
    use work.all;

entity xnoren_e is
	port(
		a_i:in	std_logic;
		b_i:in std_logic;
		en_i:in	std_logic;
		y_o: out std_logic);
end entity xnoren_e;
		


