architecture dff_a of dff_e is
	
end dff_a;
