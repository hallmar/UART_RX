library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity dff_e is
PORT(
	d_i: IN std_logic;
	clk_i: IN std_logic;
	rb_i: IN std_logic;
	en_i: IN std_logic;
	q_o: IN std_logic);
end dff_e;
